-- subtype used in design
library ieee ;
use ieee.std_logic_1164.all ;
use ieee.std_logic_arith.all ;

package cpu_types is
    type statetype is (S0, S1, S2);

    -- fix git pls
end cpu_types ;